----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:46:55 11/22/2021 
-- Design Name: 
-- Module Name:    MAIN - structural 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MAIN IS
PORT( IN1 , IN2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
          CLK , SLCT : IN STD_LOGIC;
		    OUTT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END MAIN;

ARCHITECTURE STRUCTURAL OF MAIN IS

COMPONENT REGISTE
PORT(INPUT :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	  ENABLE : IN  STD_LOGIC:='1';
     RESET : IN  STD_LOGIC:='0';
	  CLOCK : IN STD_LOGIC ;
	  OUTPUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;


COMPONENT ADDER
PORT(INPUT1 :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	  INPUT2 :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	  OUTPUT_ADD :OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;


COMPONENT MULTIPLIER
PORT(INPUT1_MUL :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	  INPUT2_MUL :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	  OUTPUT_MUL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT;


COMPONENT MULTIPLEXER
PORT(INPUT1_MUX :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	  INPUT2_MUX : IN STD_LOGIC_VECTOR(15 DOWNTO 0) ;
	  CLOCK : IN STD_LOGIC;
	  SEL : IN STD_LOGIC;
	  OUTPUT_mux : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT;

CONSTANT Z0 :STD_LOGIC:='0';
CONSTANT Z1 :STD_LOGIC:='1';
SIGNAL S1 , S2 , S3: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL S4 :STD_LOGIC_VECTOR(15 DOWNTO 0);


BEGIN

REG1:REGISTE  PORT MAP(IN1 , ENABLE=>Z1 , RESET=>Z0 , CLOCK=>CLK ,OUTPUT=>S1);

REG2:REGISTE  PORT MAP(IN2 , ENABLE=>Z1 , RESET=>Z0 , CLOCK=>CLK , OUTPUT=>S2);

ADD:ADDER     PORT MAP(S1,S2,S3);

MUL:MULTIPLIER  PORT MAP(S1,S2,S4);

MUX:MULTIPLEXER PORT MAP(S3,S4,CLK,SLCT,OUTT);


END STRUCTURAL;

